library ieee;
USE ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL; 
use IEEE.STD_LOGIC_UNSIGNED.ALL; 

ENTITY Lab7a IS
 PORT (KEY : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
 SW : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
 LEDR: OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
  LEDG: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END Lab7a;

ARCHITECTURE BEHAVIOR OF Lab7a IS 

SIGNAL CLOCK: STD_LOGIC;
SIGNAL RESET: STD_LOGIC;
SIGNAL ENTRADA: STD_LOGIC;
SIGNAL SAIDA: STD_LOGIC;
SIGNAL ESTADOP, ESTADOF: STD_LOGIC_VECTOR(8 DOWNTO 0);

COMPONENT FFD IS
	PORT (Clk, D, Clear: IN STD_LOGIC;
			Q: OUT STD_LOGIC);
END COMPONENT;
BEGIN

	LEDR(17) <= SW(17);
	ENTRADA <= SW (17);
	LEDR(8 DOWNTO 0)<=ESTADOF;
	CLOCK <= KEY(0);
	RESET <= KEY(1);
	LEDG(1 DOWNTO 0) <= KEY(1 DOWNTO 0);
	
	FF8: FFD PORT MAP(CLOCK,ESTADOP(8),RESET,ESTADOF(8));
	FF7: FFD PORT MAP(CLOCK,ESTADOP(7),RESET,ESTADOF(7));
	FF6: FFD PORT MAP(CLOCK,ESTADOP(6),RESET,ESTADOF(6));
	FF5: FFD PORT MAP(CLOCK,ESTADOP(5),RESET,ESTADOF(5));
	FF4: FFD PORT MAP(CLOCK,ESTADOP(4),RESET,ESTADOF(4));
	FF3: FFD PORT MAP(CLOCK,ESTADOP(3),RESET,ESTADOF(3));
	FF2: FFD PORT MAP(CLOCK,ESTADOP(2),RESET,ESTADOF(2));
	FF1: FFD PORT MAP(CLOCK,ESTADOP(1),RESET,ESTADOF(1));
	FF0: FFD PORT MAP(CLOCK,'1',RESET,ESTADOF(0));
	
	ESTADOP(8) <= (ESTADOF(8) AND ENTRADA) OR (ESTADOF(7) AND ENTRADA);
	ESTADOP(7) <= (ESTADOF(6) AND ENTRADA);
	ESTADOP(6) <= (ESTADOF(5) AND ENTRADA);
	ESTADOP(5) <= (NOT (ESTADOF(0)) AND ENTRADA) OR (ESTADOF(1) AND ENTRADA) OR (ESTADOF(2) AND ENTRADA) OR (ESTADOF(3) AND ENTRADA) OR (ESTADOF(4) AND ENTRADA);
	ESTADOP(4) <= (ESTADOF(4) AND NOT(ENTRADA)) OR (ESTADOF(3) AND NOT(ENTRADA));
	ESTADOP(3) <= (ESTADOF(2) AND NOT(ENTRADA));
	ESTADOP(2) <= (ESTADOF(1) AND NOT(ENTRADA));
	ESTADOP(1) <= (NOT (ESTADOF(0)) AND NOT(ENTRADA)) OR (ESTADOF(5) AND NOT(ENTRADA)) OR (ESTADOF(6) AND NOT(ENTRADA)) OR (ESTADOF(7) AND NOT(ENTRADA)) OR (ESTADOF(8) AND NOT(ENTRADA));

LEDG(4)<= ESTADOF(4) OR ESTADOF(8);

END BEHAVIOR;