library ieee;
USE ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL; 
use IEEE.STD_LOGIC_UNSIGNED.ALL; 

ENTITY Lab7b IS
 PORT (KEY : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
 SW : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
 LEDR: OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
  LEDG: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END Lab7b;

ARCHITECTURE Behavior OF Lab7b IS

SIGNAL W: STD_LOGIC;
SIGNAL CLOCK: STD_LOGIC;
SIGNAL RESET: STD_LOGIC;
SIGNAL ESTADO: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL ESTADOA: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL ESTADOB: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL ESTADOC: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL ESTADOD: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL ESTADOE: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL ESTADOF: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL ESTADOG: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL ESTADOH: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL ESTADOI: STD_LOGIC_VECTOR(8 DOWNTO 0);


TYPE State_type IS (A, B, C, D, E, F, G, H, I);
SIGNAL y_Q, y_D : State_type; 
BEGIN




W<=SW(17);
LEDR(17) <= SW(17);
CLOCK <= KEY(0);
RESET <= KEY(1);
LEDG(1 DOWNTO 0) <= KEY(1 DOWNTO 0);

	ESTADOA<="000000000";
	ESTADOB<="000000011";
	ESTADOC<="000000101";
	ESTADOD<="000001001";
	ESTADOE<="000010001";
	ESTADOF<="000100001";
	ESTADOG<="001000001";
	ESTADOH<="010000001";
	ESTADOI<="100000001";
	
PROCESS (w, y_Q)

BEGIN


	

case y_Q IS
WHEN A => IF (w = '0') THEN y_D <= B;
ELSE y_D <= F;

END IF;

WHEN B => IF (w = '0') THEN y_D <= C;
ELSE y_D <= F;

END IF;

WHEN C => IF (w = '0') THEN y_D <= D;
ELSE y_D <= F;

END IF;

WHEN D => IF (w = '0') THEN y_D <= E;
ELSE y_D <= F;

END IF;

WHEN E => IF (w = '0') THEN y_D <= E;
ELSE y_D <= F;

END IF;

WHEN F => IF (w = '0') THEN y_D <= B;
ELSE y_D <= G;

END IF;

WHEN G => IF (w = '0') THEN y_D <= B;
ELSE y_D <= H;

END IF;

WHEN H => IF (w = '0') THEN y_D <= B;
ELSE y_D <= I;


END IF;

WHEN I => IF (w = '0') THEN y_D <= B;
ELSE y_D <= I;


END IF;

END CASE;

END PROCESS; 

PROCESS (Y_Q)

BEGIN

IF(Y_Q=E OR y_Q=I) THEN
LEDG(4)<='1';
ELSE
LEDG(4)<='0';
 
 END IF;

END PROCESS;

PROCESS (Clock, RESET)
BEGIN

if (reset ='0') then
y_Q<=A;
ELSIF (rising_edge(Clock)) THEN
y_Q <= y_D;
END IF;

IF (Y_Q = A) THEN
ESTADO <= ESTADOA;
ELSIF (Y_Q = B) THEN
ESTADO <= ESTADOB;
ELSIF (Y_Q = C) THEN
ESTADO <= ESTADOC;
ELSIF (Y_Q = D) THEN
ESTADO <= ESTADOD;
ELSIF (Y_Q = E) THEN
ESTADO <= ESTADOE;
ELSIF (Y_Q = F) THEN
ESTADO <= ESTADOF;
ELSIF (Y_Q = G) THEN
ESTADO <= ESTADOG;
ELSIF (Y_Q = H) THEN
ESTADO <= ESTADOH;
ELSIF (Y_Q = I) THEN
ESTADO <= ESTADOI;
END IF;

END PROCESS;

	LEDR(17) <= SW(17);


	LEDR(8 DOWNTO 0) <= ESTADO;
	
	
	Clock <= KEY(0);
	W<=SW(17);
	RESET <= KEY(1);
	
END Behavior;

