LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY visor IS

PORT (A7: in STD_LOGIC_VECTOR(0 to 3);
		B7: out STD_LOGIC_VECTOR(0 to 6));
END visor;

		ARCHITECTURE comportamento of visor IS
		BEGIN

		B7(0 to 6) <= "0000001" WHEN A7="0000" ELSE
		"1001111" WHEN A7="0001" ELSE
		"0010010" WHEN A7="0010" ELSE
		"0000110" WHEN A7="0011" ELSE
		"1001100" WHEN A7="0100" ELSE
		"0100100" WHEN A7="0101" ELSE
		"0100000" WHEN A7="0110" ELSE
		"0001111" WHEN A7="0111" ELSE
		"0000000" WHEN A7="1000" ELSE
		"0000100" WHEN A7="1001" ELSE
		"0001000" WHEN A7="1010" ELSE
		"1100000" WHEN A7="1011" ELSE
		"0110010" WHEN A7="1100" ELSE
		"1000010" WHEN A7="1101" ELSE
		"0110000" WHEN A7="1110" ELSE
		"0111000" WHEN A7="1111" ELSE
		"1111111";
		
		END comportamento;