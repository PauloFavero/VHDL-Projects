LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Exp3e IS
PORT ( SW : IN STD_LOGIC_VECTOR (0 TO 15);
KEY: IN STD_LOGIC_vector(0 to 1);
LEDR : OUT STD_LOGIC_VECTOR(0 TO 15);
HEX0,HEX1,HEX2,HEX3,HEX4,HEX5,HEX6,HEX7: OUT STD_LOGIC_VECTOR (0 TO 6));

END Exp3e;


ARCHITECTURE BEHAVIOR OF Exp3e IS

SIGNAL FFD_VISOR4: STD_LOGIC_VECTOR(0 TO 3);
SIGNAL FFD_VISOR5: STD_LOGIC_VECTOR(0 TO 3);
SIGNAL FFD_VISOR6: STD_LOGIC_VECTOR(0 TO 3);
SIGNAL FFD_VISOR7: STD_LOGIC_VECTOR(0 TO 3);

COMPONENT FFDReset
PORT ( clk, D, rst : IN STD_LOGIC;
Q : OUT STD_LOGIC);
END COMPONENT;

COMPONENT visor
PORT (A7: in STD_LOGIC_VECTOR(0 to 3);
		B7: out STD_LOGIC_VECTOR(0 to 6));
END COMPONENT;

BEGIN 

B0: visor PORT MAP (SW(0 to 3),HEX0 (0 TO 6));
B1: visor PORT MAP (SW(4 to 7),HEX1 (0 TO 6));
B2: visor PORT MAP (SW(8 to 11),HEX2 (0 TO 6));
B3: visor PORT MAP (SW(12 to 15),HEX3 (0 TO 6));

A4_0: FFDReset PORT MAP (KEY(1),SW(0),KEY(0),FFD_VISOR4(0));
A4_1: FFDReset PORT MAP (KEY(1),SW(1),KEY(0),FFD_VISOR4(1));
A4_2: FFDReset PORT MAP (KEY(1),SW(2),KEY(0),FFD_VISOR4(2));
A4_3: FFDReset PORT MAP (KEY(1),SW(3),KEY(0),FFD_VISOR4(3));

A5_0: FFDReset PORT MAP (KEY(1),SW(4),KEY(0),FFD_VISOR5(0));
A5_1: FFDReset PORT MAP (KEY(1),SW(5),KEY(0),FFD_VISOR5(1));
A5_2: FFDReset PORT MAP (KEY(1),SW(6),KEY(0),FFD_VISOR5(2));
A5_3: FFDReset PORT MAP (KEY(1),SW(7),KEY(0),FFD_VISOR5(3));

A6_0: FFDReset PORT MAP (KEY(1),SW(8),KEY(0),FFD_VISOR6(0));
A6_1: FFDReset PORT MAP (KEY(1),SW(9),KEY(0),FFD_VISOR6(1));
A6_2: FFDReset PORT MAP (KEY(1),SW(10),KEY(0),FFD_VISOR6(2));
A6_3: FFDReset PORT MAP (KEY(1),SW(11),KEY(0),FFD_VISOR6(3));

A7_0: FFDReset PORT MAP (KEY(1),SW(12),KEY(0),FFD_VISOR7(0));
A7_1: FFDReset PORT MAP (KEY(1),SW(13),KEY(0),FFD_VISOR7(1));
A7_2: FFDReset PORT MAP (KEY(1),SW(14),KEY(0),FFD_VISOR7(2));
A7_3: FFDReset PORT MAP (KEY(1),SW(15),KEY(0),FFD_VISOR7(3));

A4: visor PORT MAP (FFD_VISOR4(0 to 3),HEX4 (0 TO 6));
A5: visor PORT MAP (FFD_VISOR5(0 to 3),HEX5 (0 TO 6));
A6: visor PORT MAP (FFD_VISOR6(0 to 3),HEX6 (0 TO 6));
A7: visor PORT MAP (FFD_VISOR7(0 to 3),HEX7 (0 TO 6));




END BEHAVIOR;