LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY visor IS

PORT (AAA7: in STD_LOGIC_VECTOR(0 to 3);
	BBB7: out STD_LOGIC_VECTOR(0 to 6));
END visor;

		ARCHITECTURE comportamento of visor IS
		BEGIN

		BBB7(0 to 6) <= "0000001" WHEN AAA7="0000" ELSE
		"1001111" WHEN AAA7="0001" ELSE
		"0010010" WHEN AAA7="0010" ELSE
		"0000110" WHEN AAA7="0011" ELSE
		"1001100" WHEN AAA7="0100" ELSE
		"0100100" WHEN AAA7="0101" ELSE
		"0100000" WHEN AAA7="0110" ELSE
		"0001111" WHEN AAA7="0111" ELSE
		"0000000" WHEN AAA7="1000" ELSE
		"0000100" WHEN AAA7="1001" ELSE
		"1111111";	
	
		
		END comportamento;